module Top_8bit(rst,clk,x0,x1,x2,x3,x4,y0,y1,y2,y3,y4);
  input rst,clk;
  input [7:0] x0,x1,x2,x3,x4;
  output [7:0] y0,y1,y2,y3,y4;
  reg [255:0] S0=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S1=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S2=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S3=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S4=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S5=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S6=256'h1243254323242343234923522342394839544352304;
  reg [255:0] S7=256'h1243254323242343234923522342394839544352304;
  Top Top1(.rst(rst),.clk(clk),.S(S0),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[0]),.y1(y1[0]),.y2(y2[0]),.y3(y3[0]),.y4(y4[0]));
  Top Top2(.rst(rst),.clk(clk),.S(S1),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[1]),.y1(y1[1]),.y2(y2[1]),.y3(y3[1]),.y4(y4[1]));
  Top Top3(.rst(rst),.clk(clk),.S(S2),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[2]),.y1(y1[2]),.y2(y2[2]),.y3(y3[2]),.y4(y4[2]));
  Top Top4(.rst(rst),.clk(clk),.S(S3),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[3]),.y1(y1[3]),.y2(y2[3]),.y3(y3[3]),.y4(y4[3]));
  Top Top5(.rst(rst),.clk(clk),.S(S4),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[4]),.y1(y1[4]),.y2(y2[4]),.y3(y3[4]),.y4(y4[4]));
  Top Top6(.rst(rst),.clk(clk),.S(S5),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[5]),.y1(y1[5]),.y2(y2[5]),.y3(y3[5]),.y4(y4[5]));
  Top Top7(.rst(rst),.clk(clk),.S(S6),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[6]),.y1(y1[6]),.y2(y2[6]),.y3(y3[6]),.y4(y4[6]));
  Top Top8(.rst(rst),.clk(clk),.S(S7),.x0(x0),.x1(x1),.x2(x2),.x3(x3),.x4(x4),.y0(y0[7]),.y1(y1[7]),.y2(y2[7]),.y3(y3[7]),.y4(y4[7]));
endmodule
